`timescale 1ns / 1ps

// n4fpga.v - Top level module for the ECE 544 Project 1
//
// Copyright Chetan Bornarkar, Portland State University, 2016
// 
// Created By:	Roy Kravitz
// Modified By: Chetan Bornarkar, Randon Stasney
// Date:		2/1/2017
// Version:		2.0
//
// Description:
// ------------
// This module provides the top level for 544 Project 1
// The module assume that a PmodOLED is plugged into the JA 
// expansion ports and that a PmodENC is plugged into the JD expansion 
// port (bottom row).  
//////////////////////////////////////////////////////////////////////
module n4fpga(
    input				clk,			// 100Mhz clock input
    input				btnC,			// center pushbutton
    input				btnU,			// UP (North) pusbhbutton
    input				btnL,			// LEFT (West) pushbutton
    input				btnD,			// DOWN (South) pushbutton  
    input				btnR,			// RIGHT (East) pushbutton
	input				btnCpuReset,	// CPU reset pushbutton
    input	[15:0]		sw,				// slide switches on Nexys 4
    output	[15:0] 		led,			// LEDs on Nexys 4   
    output              RGB1_Blue,      // RGB1 LED (LD16) 
    output              RGB1_Green,
    output              RGB1_Red,
    output              RGB2_Blue,      // RGB2 LED (LD17)
    output              RGB2_Green,
    output              RGB2_Red,
    output [7:0]        an,             // Seven Segment display
    output [6:0]        seg,
    output              dp,             // decimal point display on the seven segment 
    
    input				uart_rtl_rxd,	// USB UART Rx and Tx on Nexys 4
    output				uart_rtl_txd,	
    
	inout   [7:0]       JA,             // JA PmodOLED connector 
	                                    // both rows are used 
    inout	[7:0] 		JB,				// JB Pmod connector 
                                        // Unused. Can be used for debuggin purposes 
    inout	[7:0] 		JC,				// JC Pmod connector - debug signals
										// Can be used for debug purposes
	inout	[7:0]		JD,				// JD Pmod connector - PmodENC signals
	
	inout 			XA_N, 
	
	inout			XA_P
);

// internal variables
// Pulse Width Modulation Detecttion variables

wire				rx_sonar, tx_sonar, tx_kinect, rx_kinect;
// Clock and Reset 
wire				sysclk;              			// 100 MHz, 10 MHz
wire				sysreset_n, sysreset;					// active low reset, active high reset

// Rotary encoder 
wire				HB3_FBAR, HB3_FBAL, DIRR, ENAR, DIRL, ENAL;
wire 	[3:0]		Arduino_Enc;

// GPIO pins 
wire	[31:0]	    gpio_in;				// embsys GPIO input port
wire	[31:0]	    gpio_out;				// embsys GPIO output port

// OLED pins 
wire 				pmodoledrgb_out_pin1_i, pmodoledrgb_out_pin1_io, pmodoledrgb_out_pin1_o, pmodoledrgb_out_pin1_t; 
wire 				pmodoledrgb_out_pin2_i, pmodoledrgb_out_pin2_io, pmodoledrgb_out_pin2_o, pmodoledrgb_out_pin2_t; 
wire 				pmodoledrgb_out_pin3_i, pmodoledrgb_out_pin3_io, pmodoledrgb_out_pin3_o, pmodoledrgb_out_pin3_t; 
wire 				pmodoledrgb_out_pin4_i, pmodoledrgb_out_pin4_io, pmodoledrgb_out_pin4_o, pmodoledrgb_out_pin4_t; 
wire 				pmodoledrgb_out_pin7_i, pmodoledrgb_out_pin7_io, pmodoledrgb_out_pin7_o, pmodoledrgb_out_pin7_t; 
wire 				pmodoledrgb_out_pin8_i, pmodoledrgb_out_pin8_io, pmodoledrgb_out_pin8_o, pmodoledrgb_out_pin8_t; 
wire 				pmodoledrgb_out_pin9_i, pmodoledrgb_out_pin9_io, pmodoledrgb_out_pin9_o, pmodoledrgb_out_pin9_t; 
wire 				pmodoledrgb_out_pin10_i, pmodoledrgb_out_pin10_io, pmodoledrgb_out_pin10_o, pmodoledrgb_out_pin10_t;

wire 				pmodbt_out_pin1_i, pmodbt_out_pin1_io, pmodbt_out_pin1_o, pmodbt_out_pin1_t; 
wire 				pmodbt_out_pin2_i, pmodbt_out_pin2_io, pmodbt_out_pin2_o, pmodbt_out_pin2_t; 
wire 				pmodbt_out_pin3_i, pmodbt_out_pin3_io, pmodbt_out_pin3_o, pmodbt_out_pin3_t; 
wire 				pmodbt_out_pin4_i, pmodbt_out_pin4_io, pmodbt_out_pin4_o, pmodbt_out_pin4_t; 
wire 				pmodbt_out_pin7_i, pmodbt_out_pin7_io, pmodbt_out_pin7_o, pmodbt_out_pin7_t; 
wire 				pmodbt_out_pin8_i, pmodbt_out_pin8_io, pmodbt_out_pin8_o, pmodbt_out_pin8_t; 
wire 				pmodbt_out_pin9_i, pmodbt_out_pin9_io, pmodbt_out_pin9_o, pmodbt_out_pin9_t; 
wire 				pmodbt_out_pin10_i, pmodbt_out_pin10_io, pmodbt_out_pin10_o, pmodbt_out_pin10_t;

// RGB LED 
wire                w_RGB1_Red, w_RGB1_Blue, w_RGB1_Green;

// PWMDET RGB
wire 				[6:0] PW_Red;			// Red duty cycle as 7 bit value
wire 				[6:0] PW_Green;			// Green duty cycle as 7 bit value
wire 				[6:0] PW_Blue;			// Blue duty cycle as 7 bit value
// LED pins 
wire    [15:0]      led_int;                // Nexys4IO drives these outputs



assign sysclk = clk;
// connect driving wires back through gpio for SW PWMDet	
assign w_RGB1_Red = RGB1_Red;
assign w_RGB1_Blue = RGB1_Blue;
assign w_RGB1_Green = RGB1_Green;

// connect the HW PWMDet to be returned to microblaze
//assign PW_Blue = blue_test[6:0];
//assign PW_Red = red_test[6:0];
//assign PW_Green = green_test[6:0];

assign Arduino_Enc = JC [3:0];
assign gpio_in = {28'b0, Arduino_Enc};

// Drive the leds from the signal generated by the microblaze 
assign led = led_int;                   // LEDs are driven by led

// make the connections
// system-wide signals
assign sysreset_n = btnCpuReset;		// The CPU reset pushbutton is asserted low.  The other pushbuttons are asserted high
										// but the microblaze for Nexys 4 expects reset to be asserted low
assign sysreset = ~sysreset_n;			// Generate a reset signal that is asserted high for any logic blocks expecting it.

// Pmod OLED connections 
assign JB[0] = pmodoledrgb_out_pin1_io;
assign JB[1] = pmodoledrgb_out_pin2_io;
assign JB[2] = pmodoledrgb_out_pin3_io;
assign JB[3] = pmodoledrgb_out_pin4_io;
assign JB[4] = pmodoledrgb_out_pin7_io;
assign JB[5] = pmodoledrgb_out_pin8_io;
assign JB[6] = pmodoledrgb_out_pin9_io;
assign JB[7] = pmodoledrgb_out_pin10_io;
//rx_sonar, tx_kinect;
// JB Connector connections can be used for debug purposes
//assign tx_kinect = JA[0];
//assign JA[1] = rx_kinect;

//assign tx_sonar = JA[5];
//assign JA[6] = rx_sonar;

//ssign JD[1] = pmodbt_out_pin2_io;
assign JA[0] = pmodbt_out_pin1_io;
assign JA[1] = pmodbt_out_pin2_io;
assign JA[2] = pmodbt_out_pin3_io;
assign JA[3] = pmodbt_out_pin4_io;
assign JA[4] = pmodbt_out_pin7_io;
assign JA[5] = pmodbt_out_pin8_io;
assign JA[6] = pmodbt_out_pin9_io;
assign JA[7] = pmodbt_out_pin10_io;

// JC Connector pins can be used for debug purposes 
//assign JC[3:0] = 4'h0; 
assign JD[4] = DIRL;
assign JD[5] = ENAL;
assign HB3_FBAR = JD[6];
assign JD[7] = 1'b0;
assign JC[4] = DIRR;
assign JC[5] = ENAR;
assign HB3_FBAR = JC[6];
assign  JC[7] = 1'b0;
//assign DIR = 1'b0;
//assign ENA = RGB1_Blue;
//HB3_FBA, HB3_FBB, DIR, ENA
// PmodENC signals
// JD - bottom row only
// Pins are assigned such that turning the knob to the right
// causes the rotary count to increment.
//assign rotary_a = JA[5];
//assign rotary_b = JA[4];
//assign rotary_press = JA[6];
//assign rotary_sw = JA[7];
/*
// simple block for hardware detection
always @ (posedge detclk)
begin	// default assigments to avoid latches
		blue_test <= blue_test;								
		blue_test_count <= blue_test_count;
		red_test <= red_test;
		red_test_count <= red_test_count;
		green_test <= green_test;
		green_test_count <= green_test_count;
		
	if (time_base == 0)										// 6,400,000 count reaches zero
		begin
		time_base <= 23'b110_0001_1010_1000_0000_0000;		// reset count
		blue_test_count <= 0;								// reset high counts
		blue_test <= blue_test_count/64000;					// calculate detected blue duty cycle
		red_test_count <= 0;								// reset high counts
		red_test <= red_test_count/64000;					// calculate detected red duty cycle
		green_test_count <= 0;								// reset high counts
		green_test <= green_test_count/64000;				// // calculate detected green duty cycle
		end
	else													// otherwise
		begin
		time_base <= time_base - 1;							// decrement counter
		if (RGB1_Blue == 1)
		blue_test_count <= blue_test_count + 1;				// if signal high increment count
		if (HB3_FBA == 1)
		red_test_count <= red_test_count + 1;				// if signal high increment count
//if (HB3_FBA == 1)
		green_test_count <= green_test_count + 1;			// if signal high increment count
		end
end
*/
// instantiate the embedded system
design_1 Design_1
       (// PMOD OLED pins 
        .PmodOLEDrgb_out_pin10_i(pmodoledrgb_out_pin10_i),
	    .PmodOLEDrgb_out_pin10_o(pmodoledrgb_out_pin10_o),
	    .PmodOLEDrgb_out_pin10_t(pmodoledrgb_out_pin10_t),
	    .PmodOLEDrgb_out_pin1_i(pmodoledrgb_out_pin1_i),
	    .PmodOLEDrgb_out_pin1_o(pmodoledrgb_out_pin1_o),
	    .PmodOLEDrgb_out_pin1_t(pmodoledrgb_out_pin1_t),
	    .PmodOLEDrgb_out_pin2_i(pmodoledrgb_out_pin2_i),
	    .PmodOLEDrgb_out_pin2_o(pmodoledrgb_out_pin2_o),
	    .PmodOLEDrgb_out_pin2_t(pmodoledrgb_out_pin2_t),
	    .PmodOLEDrgb_out_pin3_i(pmodoledrgb_out_pin3_i),
	    .PmodOLEDrgb_out_pin3_o(pmodoledrgb_out_pin3_o),
	    .PmodOLEDrgb_out_pin3_t(pmodoledrgb_out_pin3_t),
	    .PmodOLEDrgb_out_pin4_i(pmodoledrgb_out_pin4_i),
	    .PmodOLEDrgb_out_pin4_o(pmodoledrgb_out_pin4_o),
	    .PmodOLEDrgb_out_pin4_t(pmodoledrgb_out_pin4_t),
	    .PmodOLEDrgb_out_pin7_i(pmodoledrgb_out_pin7_i),
	    .PmodOLEDrgb_out_pin7_o(pmodoledrgb_out_pin7_o),
	    .PmodOLEDrgb_out_pin7_t(pmodoledrgb_out_pin7_t),
	    .PmodOLEDrgb_out_pin8_i(pmodoledrgb_out_pin8_i),
	    .PmodOLEDrgb_out_pin8_o(pmodoledrgb_out_pin8_o),
	    .PmodOLEDrgb_out_pin8_t(pmodoledrgb_out_pin8_t),
	    .PmodOLEDrgb_out_pin9_i(pmodoledrgb_out_pin9_i),
	    .PmodOLEDrgb_out_pin9_o(pmodoledrgb_out_pin9_o),
	    .PmodOLEDrgb_out_pin9_t(pmodoledrgb_out_pin9_t),
		
        .Pmod_out_pin10_i(pmodbt_out_pin10_i),
	    .Pmod_out_pin10_o(pmodbt_out_pin10_o),
	    .Pmod_out_pin10_t(pmodbt_out_pin10_t),
	    .Pmod_out_pin1_i(pmodbt_out_pin1_i),
	    .Pmod_out_pin1_o(pmodbt_out_pin1_o),
	    .Pmod_out_pin1_t(pmodbt_out_pin1_t),
	    .Pmod_out_pin2_i(pmodbt_out_pin2_i),
	    .Pmod_out_pin2_o(pmodbt_out_pin2_o),
	    .Pmod_out_pin2_t(pmodbt_out_pin2_t),
	    .Pmod_out_pin3_i(pmodbt_out_pin3_i),
	    .Pmod_out_pin3_o(pmodbt_out_pin3_o),
	    .Pmod_out_pin3_t(pmodbt_out_pin3_t),
	    .Pmod_out_pin4_i(pmodbt_out_pin4_i),
	    .Pmod_out_pin4_o(pmodbt_out_pin4_o),
	    .Pmod_out_pin4_t(pmodbt_out_pin4_t),
	    .Pmod_out_pin7_i(pmodbt_out_pin7_i),
	    .Pmod_out_pin7_o(pmodbt_out_pin7_o),
	    .Pmod_out_pin7_t(pmodbt_out_pin7_t),
	    .Pmod_out_pin8_i(pmodbt_out_pin8_i),
	    .Pmod_out_pin8_o(pmodbt_out_pin8_o),
	    .Pmod_out_pin8_t(pmodbt_out_pin8_t),
	    .Pmod_out_pin9_i(pmodbt_out_pin9_i),
	    .Pmod_out_pin9_o(pmodbt_out_pin9_o),
	    .Pmod_out_pin9_t(pmodbt_out_pin9_t),

	    // GPIO pins 
  //  gpio_0_GPIO2_tri_i,
   //     gpio_0_GPIO_tri_o,
        .gpio_0_GPIO_tri_i(gpio_in),
        .gpio_0_GPIO2_tri_o(gpio_out),
        // Pmod Rotary Encoder
	   // .pmodENC_A(rotary_a),
       // .pmodENC_B(rotary_b),
       // .pmodENC_btn(rotary_press),
       // .pmodENC_sw(rotary_sw),
        // RGB1/2 Led's 
        .RGB1_Blue(RGB1_Blue),
        .RGB1_Green(RGB1_Green),
        .RGB1_Red(RGB1_Red),
        .RGB2_Blue(RGB2_Blue),
        .RGB2_Green(RGB2_Green),
        .RGB2_Red(RGB2_Red),
        // Seven Segment Display anode control  
        .an(an),
        .dp(dp),
        .led(led_int),
        .seg(seg),
        // Push buttons and switches  
        .btnC(btnC),
        .btnD(btnD),
        .btnL(btnL),
        .btnR(btnR),
        .btnU(btnU),
        .sw(sw),
        // reset and clock 
        .sysreset_n(sysreset_n),
        .sysclk(sysclk),
        // UART pins 
		.Vaux3_v_n(XA_N),
		.Vaux3_v_p(XA_P),
		
		
    //.uart_rtl_0_rxd(tx_kinect),
    //.uart_rtl_0_txd(rx_kinect),
    //.uart_rtl_1_rxd(tx_sonar),
    //.uart_rtl_1_txd(rx_sonar),
     
        .uart_rtl_rxd(uart_rtl_rxd),
        .uart_rtl_txd(uart_rtl_txd),
		// HB3
		.ENABLE(ENAL),
		.DIRECTION(DIRR),
		.SA(HB3_FBAR),
		.SB(1'b1),
		.ENABLE_1(ENAR),
		.DIRECTION_1(DIRL),
		.SA_1(HB3_FBAL),


		.SB_1(1'b1)
);
     
// Tristate buffers for the pmodOLEDrgb pins
// generated by PMOD bridge component.  Many
// of these signals are not tri-state.
IOBUF pmodbt_out_pin1_iobuf
(
    .I(pmodbt_out_pin1_o),
    .IO(pmodbt_out_pin1_io),
    .O(pmodbt_out_pin1_i),
    .T(pmodbt_out_pin1_t)
);

IOBUF pmodbt_out_pin2_iobuf
(
    .I(pmodbt_out_pin2_o),
    .IO(pmodbt_out_pin2_io),
    .O(pmodbt_out_pin2_i),
    .T(pmodbt_out_pin2_t)
);

IOBUF pmodbt_out_pin3_iobuf
(
    .I(pmodbt_out_pin3_o),
    .IO(pmodbt_out_pin3_io),
    .O(pmodbt_out_pin3_i),
    .T(pmodbt_out_pin3_t)
);

IOBUF pmodbt_out_pin4_iobuf
(
    .I(pmodbt_out_pin4_o),
    .IO(pmodbt_out_pin4_io),
    .O(pmodbt_out_pin4_i),
    .T(pmodbt_out_pin4_t)
);

IOBUF pmodbt_out_pin7_iobuf
(
    .I(pmodbt_out_pin7_o),
    .IO(pmodbt_out_pin7_io),
    .O(pmodbt_out_pin7_i),
    .T(pmodbt_out_pin7_t)
);

IOBUF pmodbt_out_pin8_iobuf
(
    .I(pmodbt_out_pin8_o),
    .IO(pmodbt_out_pin8_io),
    .O(pmodbt_out_pin8_i),
    .T(pmodbt_out_pin8_t)
);

IOBUF pmodbt_out_pin9_iobuf
(
    .I(pmodbt_out_pin9_o),
    .IO(pmodbt_out_pin9_io),
    .O(pmodbt_out_pin9_i),
    .T(pmodbt_out_pin9_t)
);

IOBUF pmodbt_out_pin10_iobuf
(
    .I(pmodbt_out_pin10_o),
    .IO(pmodbt_out_pin10_io),
    .O(pmodbt_out_pin10_i),
    .T(pmodbt_out_pin10_t)
);

IOBUF pmodoledrgb_out_pin1_iobuf
(
    .I(pmodoledrgb_out_pin1_o),
    .IO(pmodoledrgb_out_pin1_io),
    .O(pmodoledrgb_out_pin1_i),
    .T(pmodoledrgb_out_pin1_t)
);

IOBUF pmodoledrgb_out_pin2_iobuf
(
    .I(pmodoledrgb_out_pin2_o),
    .IO(pmodoledrgb_out_pin2_io),
    .O(pmodoledrgb_out_pin2_i),
    .T(pmodoledrgb_out_pin2_t)
);

IOBUF pmodoledrgb_out_pin3_iobuf
(
    .I(pmodoledrgb_out_pin3_o),
    .IO(pmodoledrgb_out_pin3_io),
    .O(pmodoledrgb_out_pin3_i),
    .T(pmodoledrgb_out_pin3_t)
);

IOBUF pmodoledrgb_out_pin4_iobuf
(
    .I(pmodoledrgb_out_pin4_o),
    .IO(pmodoledrgb_out_pin4_io),
    .O(pmodoledrgb_out_pin4_i),
    .T(pmodoledrgb_out_pin4_t)
);

IOBUF pmodoledrgb_out_pin7_iobuf
(
    .I(pmodoledrgb_out_pin7_o),
    .IO(pmodoledrgb_out_pin7_io),
    .O(pmodoledrgb_out_pin7_i),
    .T(pmodoledrgb_out_pin7_t)
);

IOBUF pmodoledrgb_out_pin8_iobuf
(
    .I(pmodoledrgb_out_pin8_o),
    .IO(pmodoledrgb_out_pin8_io),
    .O(pmodoledrgb_out_pin8_i),
    .T(pmodoledrgb_out_pin8_t)
);

IOBUF pmodoledrgb_out_pin9_iobuf
(
    .I(pmodoledrgb_out_pin9_o),
    .IO(pmodoledrgb_out_pin9_io),
    .O(pmodoledrgb_out_pin9_i),
    .T(pmodoledrgb_out_pin9_t)
);

IOBUF pmodoledrgb_out_pin10_iobuf
(
    .I(pmodoledrgb_out_pin10_o),
    .IO(pmodoledrgb_out_pin10_io),
    .O(pmodoledrgb_out_pin10_i),
    .T(pmodoledrgb_out_pin10_t)
);


endmodule