`timescale 1ns / 1ps

// n4fpga.v - Top level module for the ECE 544 Getting Started project
//
// Copyright Chetan Bornarkar, Portland State University, 2016
// 
// Created By:	Roy Kravitz
// Modified By: Chetan Bornarkar
// Date:		23-December-2016
// Version:		1.0
//
// Description:
// ------------
// This module provides the top level for the Getting Started hardware.
// The module assume that a PmodOLED is plugged into the JA 
// expansion ports and that a PmodENC is plugged into the JD expansion 
// port (bottom row).  
//////////////////////////////////////////////////////////////////////
module n4fpga(
    input				clk,			// 100Mhz clock input
    input				btnC,			// center pushbutton
    input				btnU,			// UP (North) pusbhbutton
    input				btnL,			// LEFT (West) pushbutton
    input				btnD,			// DOWN (South) pushbutton  - used for system reset
    input				btnR,			// RIGHT (East) pushbutton
	input				btnCpuReset,	// CPU reset pushbutton
    input	[15:0]		sw,				// slide switches on Nexys 4
    output	[15:0] 		led,			// LEDs on Nexys 4   
    output              RGB1_Blue,      // RGB1 LED (LD16) 
    output              RGB1_Green,
    output              RGB1_Red,
    output              RGB2_Blue,      // RGB2 LED (LD17)
    output              RGB2_Green,
    output              RGB2_Red,
    output [7:0]        an,             // Seven Segment display
    output [6:0]        seg,
    output              dp,             // decimal point display on the seven segment 
    
    input				uart_rtl_rxd,	// USB UART Rx and Tx on Nexys 4
    output				uart_rtl_txd,	
    
	inout   [7:0]       JA,             // JA PmodOLED connector 
	                                    // both rows are used 
    inout	[7:0] 		JB,				// JB Pmod connector 
                                        // Unused. Can be used for debuggin purposes 
    output	[7:0] 		JC,				// JC Pmod connector - debug signals
										// Can be used for debug purposes
	input	[7:0]		JD,				// JD Pmod connector - PmodENC signals
    input               vauxn3,         //input for ADC
    input               vauxp3          //input for ADC
);

// internal variables
// Clock and Reset 
wire				sysclk;             // 
wire				sysreset_n, sysreset;

wire                uart_rx;

// Rotary encoder 
wire				rotary_a, rotary_b, rotary_press, rotary_sw;

// GPIO pins 
wire	[7:0]	    gpio_in;				// embsys GPIO input port
wire	[7:0]	    gpio_out;				// embsys GPIO output port

// OLED pins 
wire 				pmodoledrgb_out_pin1_i, pmodoledrgb_out_pin1_io, pmodoledrgb_out_pin1_o, pmodoledrgb_out_pin1_t; 
wire 				pmodoledrgb_out_pin2_i, pmodoledrgb_out_pin2_io, pmodoledrgb_out_pin2_o, pmodoledrgb_out_pin2_t; 
wire 				pmodoledrgb_out_pin3_i, pmodoledrgb_out_pin3_io, pmodoledrgb_out_pin3_o, pmodoledrgb_out_pin3_t; 
wire 				pmodoledrgb_out_pin4_i, pmodoledrgb_out_pin4_io, pmodoledrgb_out_pin4_o, pmodoledrgb_out_pin4_t; 
wire 				pmodoledrgb_out_pin7_i, pmodoledrgb_out_pin7_io, pmodoledrgb_out_pin7_o, pmodoledrgb_out_pin7_t; 
wire 				pmodoledrgb_out_pin8_i, pmodoledrgb_out_pin8_io, pmodoledrgb_out_pin8_o, pmodoledrgb_out_pin8_t; 
wire 				pmodoledrgb_out_pin9_i, pmodoledrgb_out_pin9_io, pmodoledrgb_out_pin9_o, pmodoledrgb_out_pin9_t; 
wire 				pmodoledrgb_out_pin10_i, pmodoledrgb_out_pin10_io, pmodoledrgb_out_pin10_o, pmodoledrgb_out_pin10_t;

//Bluetooth Pins
wire 				BT_out_pin1_i, BT_out_pin1_io, BT_out_pin1_o, BT_out_pin1_t; 
wire 				BT_out_pin2_i, BT_out_pin2_io, BT_out_pin2_o, BT_out_pin2_t; 
wire 				BT_out_pin3_i, BT_out_pin3_io, BT_out_pin3_o, BT_out_pin3_t; 
wire 				BT_out_pin4_i, BT_out_pin4_io, BT_out_pin4_o, BT_out_pin4_t; 
wire 				BT_out_pin7_i, BT_out_pin7_io, BT_out_pin7_o, BT_out_pin7_t; 
wire 				BT_out_pin8_i, BT_out_pin8_io, BT_out_pin8_o, BT_out_pin8_t; 
wire 				BT_out_pin9_i, BT_out_pin9_io, BT_out_pin9_o, BT_out_pin9_t; 
wire 				BT_out_pin10_i, BT_out_pin10_io, BT_out_pin10_o, BT_out_pin10_t;

// RGB LED 
wire                w_RGB1_Red, w_RGB1_Blue, w_RGB1_Green;

// LED pins 
wire    [15:0]      led_int;                // Nexys4IO drives these outputs

//motor control signals
wire                motor_pwm_out;
wire                motor_pwm_out_1;
wire                motor_sw;
wire                motor_sw_1;

// make the connections to the GPIO port.  Most of the bits are unused in the Getting
// Started project but GPIO's provide a convenient way to get the inputs and
// outputs from logic you create to and from the Microblaze.  For example,
// you may decide that using an axi_gpio peripheral is a good way to interface
// your hardware pulse-width detect logic with the Microblaze.  Our application
// is simple.
// Wrap the RGB led output back to the application program for software pulse-width detect
assign gpio_in = {5'b00000, w_RGB1_Red, w_RGB1_Blue, w_RGB1_Green};

// Drive the leds from the signal generated by the microblaze 
assign led = led_int;                   // LEDs are driven by led

// make the connections
// system-wide signals
assign sysclk = clk;
assign sysreset_n = btnCpuReset;		// The CPU reset pushbutton is asserted low.  The other pushbuttons are asserted high
										// but the microblaze for Nexys 4 expects reset to be asserted low
assign sysreset = ~sysreset_n;			// Generate a reset signal that is asserted high for any logic blocks expecting it.

// Pmod OLED connections 
assign JA[0] = pmodoledrgb_out_pin1_io;
assign JA[1] = pmodoledrgb_out_pin2_io;
assign JA[2] = pmodoledrgb_out_pin3_io;
assign JA[3] = pmodoledrgb_out_pin4_io;
assign JA[4] = pmodoledrgb_out_pin7_io;
assign JA[5] = pmodoledrgb_out_pin8_io;
assign JA[6] = pmodoledrgb_out_pin9_io;
assign JA[7] = pmodoledrgb_out_pin10_io;

// Bluetooth connections 
assign JB[0] = BT_out_pin1_io;
assign JB[1] = BT_out_pin2_io;
assign JB[2] = BT_out_pin3_io;
assign JB[3] = BT_out_pin4_io;
assign JB[4] = BT_out_pin7_io;
assign JB[5] = BT_out_pin8_io;
assign JB[6] = BT_out_pin9_io;
assign JB[7] = BT_out_pin10_io;

//motor control assignments
assign JC[0] = motor_pwm_out;
assign uart_rx = JC[1];
assign JC[3] = motor_pwm_out_1;


// instantiate the embedded system
embsys EMBSYS
       (// PMOD OLED pins 
        .PmodOLEDrgb_out_pin10_i(pmodoledrgb_out_pin10_i),
	    .PmodOLEDrgb_out_pin10_o(pmodoledrgb_out_pin10_o),
	    .PmodOLEDrgb_out_pin10_t(pmodoledrgb_out_pin10_t),
	    .PmodOLEDrgb_out_pin1_i(pmodoledrgb_out_pin1_i),
	    .PmodOLEDrgb_out_pin1_o(pmodoledrgb_out_pin1_o),
	    .PmodOLEDrgb_out_pin1_t(pmodoledrgb_out_pin1_t),
	    .PmodOLEDrgb_out_pin2_i(pmodoledrgb_out_pin2_i),
	    .PmodOLEDrgb_out_pin2_o(pmodoledrgb_out_pin2_o),
	    .PmodOLEDrgb_out_pin2_t(pmodoledrgb_out_pin2_t),
	    .PmodOLEDrgb_out_pin3_i(pmodoledrgb_out_pin3_i),
	    .PmodOLEDrgb_out_pin3_o(pmodoledrgb_out_pin3_o),
	    .PmodOLEDrgb_out_pin3_t(pmodoledrgb_out_pin3_t),
	    .PmodOLEDrgb_out_pin4_i(pmodoledrgb_out_pin4_i),
	    .PmodOLEDrgb_out_pin4_o(pmodoledrgb_out_pin4_o),
	    .PmodOLEDrgb_out_pin4_t(pmodoledrgb_out_pin4_t),
	    .PmodOLEDrgb_out_pin7_i(pmodoledrgb_out_pin7_i),
	    .PmodOLEDrgb_out_pin7_o(pmodoledrgb_out_pin7_o),
	    .PmodOLEDrgb_out_pin7_t(pmodoledrgb_out_pin7_t),
	    .PmodOLEDrgb_out_pin8_i(pmodoledrgb_out_pin8_i),
	    .PmodOLEDrgb_out_pin8_o(pmodoledrgb_out_pin8_o),
	    .PmodOLEDrgb_out_pin8_t(pmodoledrgb_out_pin8_t),
	    .PmodOLEDrgb_out_pin9_i(pmodoledrgb_out_pin9_i),
	    .PmodOLEDrgb_out_pin9_o(pmodoledrgb_out_pin9_o),
	    .PmodOLEDrgb_out_pin9_t(pmodoledrgb_out_pin9_t),
        //BT Pins
        .BT_out_pin10_i(BT_out_pin10_i),
        .BT_out_pin10_o(BT_out_pin10_o),
        .BT_out_pin10_t(BT_out_pin10_t),
        .BT_out_pin1_i(BT_out_pin1_i),
        .BT_out_pin1_o(BT_out_pin1_o),
        .BT_out_pin1_t(BT_out_pin1_t),
        .BT_out_pin2_i(BT_out_pin2_i),
        .BT_out_pin2_o(BT_out_pin2_o),
        .BT_out_pin2_t(BT_out_pin2_t),
        .BT_out_pin3_i(BT_out_pin3_i),
        .BT_out_pin3_o(BT_out_pin3_o),
        .BT_out_pin3_t(BT_out_pin3_t),
        .BT_out_pin4_i(BT_out_pin4_i),
        .BT_out_pin4_o(BT_out_pin4_o),
        .BT_out_pin4_t(BT_out_pin4_t),
        .BT_out_pin7_i(BT_out_pin7_i),
        .BT_out_pin7_o(BT_out_pin7_o),
        .BT_out_pin7_t(BT_out_pin7_t),
        .BT_out_pin8_i(BT_out_pin8_i),
        .BT_out_pin8_o(BT_out_pin8_o),
        .BT_out_pin8_t(BT_out_pin8_t),
        .BT_out_pin9_i(BT_out_pin9_i),
        .BT_out_pin9_o(BT_out_pin9_o),
        .BT_out_pin9_t(BT_out_pin9_t),
	    // GPIO pins 
//        .gpio_0_GPIO_tri_i(gpio_in),
//        .gpio_0_GPIO2_tri_o(gpio_out),
        // Pmod Rotary Encoder
//	    .pmodENC_A(rotary_a),
//        .pmodENC_B(rotary_b),
//        .pmodENC_btn(rotary_press),
//        .pmodENC_sw(rotary_sw),
        // RGB1/2 Led's 
        .RGB1_Blue(RGB1_Blue),
        .RGB1_Green(RGB1_Green),
        .RGB1_Red(RGB1_Red),
        .RGB2_Blue(RGB2_Blue),
        .RGB2_Green(RGB2_Green),
        .RGB2_Red(RGB2_Red),
        // Seven Segment Display anode control  
        .an(an),
        .dp(dp),
        .led(led_int),
        .seg(seg),
        // Push buttons and switches  
        .btnC(btnC),
        .btnD(btnD),
        .btnL(btnL),
        .btnR(btnR),
        .btnU(btnU),
        .sw(sw),
        // reset and clock 
        .sysreset_n(sysreset_n),
        .sysclk(sysclk),
        // UART pins 
        .uart_rtl_rxd(uart_rtl_rxd),
        .uart_rtl_txd(uart_rtl_txd),
        //uart for ultrasonic sensor
        .uart_rx(uart_rx),
        //Motor Control Pins
        .motor_pwm_out(motor_pwm_out),
        .motor_pwm_out_1(motor_pwm_out_1),
        .motor_sw(sw[15]),
        .motor_sw_1(sw[14]),
        .vauxn3(vauxn3),
        .vauxp3(vauxp3));
        
// Tristate buffers for the pmodOLEDrgb pins
// generated by PMOD bridge component.  Many
// of these signals are not tri-state.
IOBUF pmodoledrgb_out_pin1_iobuf
(
    .I(pmodoledrgb_out_pin1_o),
    .IO(pmodoledrgb_out_pin1_io),
    .O(pmodoledrgb_out_pin1_i),
    .T(pmodoledrgb_out_pin1_t)
);

IOBUF pmodoledrgb_out_pin2_iobuf
(
    .I(pmodoledrgb_out_pin2_o),
    .IO(pmodoledrgb_out_pin2_io),
    .O(pmodoledrgb_out_pin2_i),
    .T(pmodoledrgb_out_pin2_t)
);

IOBUF pmodoledrgb_out_pin3_iobuf
(
    .I(pmodoledrgb_out_pin3_o),
    .IO(pmodoledrgb_out_pin3_io),
    .O(pmodoledrgb_out_pin3_i),
    .T(pmodoledrgb_out_pin3_t)
);

IOBUF pmodoledrgb_out_pin4_iobuf
(
    .I(pmodoledrgb_out_pin4_o),
    .IO(pmodoledrgb_out_pin4_io),
    .O(pmodoledrgb_out_pin4_i),
    .T(pmodoledrgb_out_pin4_t)
);

IOBUF pmodoledrgb_out_pin7_iobuf
(
    .I(pmodoledrgb_out_pin7_o),
    .IO(pmodoledrgb_out_pin7_io),
    .O(pmodoledrgb_out_pin7_i),
    .T(pmodoledrgb_out_pin7_t)
);

IOBUF pmodoledrgb_out_pin8_iobuf
(
    .I(pmodoledrgb_out_pin8_o),
    .IO(pmodoledrgb_out_pin8_io),
    .O(pmodoledrgb_out_pin8_i),
    .T(pmodoledrgb_out_pin8_t)
);

IOBUF pmodoledrgb_out_pin9_iobuf
(
    .I(pmodoledrgb_out_pin9_o),
    .IO(pmodoledrgb_out_pin9_io),
    .O(pmodoledrgb_out_pin9_i),
    .T(pmodoledrgb_out_pin9_t)
);

IOBUF pmodoledrgb_out_pin10_iobuf
(
    .I(pmodoledrgb_out_pin10_o),
    .IO(pmodoledrgb_out_pin10_io),
    .O(pmodoledrgb_out_pin10_i),
    .T(pmodoledrgb_out_pin10_t)
);


// Tristate buffers for the BT module pins
IOBUF BT_out_pin1_iobuf
(
    .I(BT_out_pin1_o),
    .IO(BT_out_pin1_io),
    .O(BT_out_pin1_i),
    .T(BT_out_pin1_t)
);

IOBUF BT_out_pin2_iobuf
(
    .I(BT_out_pin2_o),
    .IO(BT_out_pin2_io),
    .O(BT_out_pin2_i),
    .T(BT_out_pin2_t)
);

IOBUF BT_out_pin3_iobuf
(
    .I(BT_out_pin3_o),
    .IO(BT_out_pin3_io),
    .O(BT_out_pin3_i),
    .T(BT_out_pin3_t)
);

IOBUF BT_out_pin4_iobuf
(
    .I(BT_out_pin4_o),
    .IO(BT_out_pin4_io),
    .O(BT_out_pin4_i),
    .T(BT_out_pin4_t)
);

IOBUF BT_out_pin7_iobuf
(
    .I(BT_out_pin7_o),
    .IO(BT_out_pin7_io),
    .O(BT_out_pin7_i),
    .T(BT_out_pin7_t)
);

IOBUF BT_out_pin8_iobuf
(
    .I(BT_out_pin8_o),
    .IO(BT_out_pin8_io),
    .O(BT_out_pin8_i),
    .T(BT_out_pin8_t)
);

IOBUF BT_out_pin9_iobuf
(
    .I(BT_out_pin9_o),
    .IO(BT_out_pin9_io),
    .O(BT_out_pin9_i),
    .T(BT_out_pin9_t)
);

IOBUF BT_out_pin10_iobuf
(
    .I(BT_out_pin10_o),
    .IO(BT_out_pin10_io),
    .O(BT_out_pin10_i),
    .T(BT_out_pin10_t)
);


endmodule

